//-- Megaherzios  MHz
`define F_50MHz 2
`define F_10MHz 10
`define F_1MHz 100
    
//-- Hertzios (Hz)
`define F_2Hz   50_000_000
`define F_1Hz   100_000_000
