module Nand(a,b, out);
  input a;
  input b;
  output out;
  nand(out,a,b);
endmodule

