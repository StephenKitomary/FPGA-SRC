// clk_in 100MHz 
`define B230400 434
`define B115200 868
`define B9600	10417
